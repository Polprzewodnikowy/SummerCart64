`define VERSION         "a"

`define BANK_INVALID    4'd0
`define BANK_SDRAM      4'd1
`define BANK_CART       4'd2
`define BANK_EEPROM     4'd3
`define BANK_SD         4'd4
